module halfadd(input wire a, b, output wire sum, cout);

 -----------------
------------------  
endmodule
