module fulladd(input wire a, b, cin, output wire sum, cout);
wire [4:0] t;

    xor2 x0(a,b,t[0]);
    xor2 x1(t[0],cin,sum);

    and2 a0(a,b,t[1]);
    and2 a1(a,cin,t[2]);
    and2 a2(b,cin,t[3]);

    or2 o0(t[1],t[2],t[4]);
    or2 o1(t[4],t[3],cout);
endmodule
